`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:07:35 12/23/2010 
// Design Name: 
// Module Name:    prom_DMH 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module prom_DMH(

input wire [3:0] addr,
input wire [7:0] key_code,
output reg [0:31] M
    );

reg [0:31] rom_A [0:15];
reg [0:31] rom_B [0:15];
reg [0:31] rom_C [0:15];
reg [0:31] rom_D [0:15];
reg [0:31] rom_E [0:15];
reg [0:31] rom_F [0:15];
reg [0:31] rom_G [0:15];
reg [0:31] rom_H [0:15];
reg [0:31] rom_I [0:15];
reg [0:31] rom_J [0:15];
reg [0:31] rom_K [0:15];
reg [0:31] rom_L [0:15];
reg [0:31] rom_M [0:15];
reg [0:31] rom_N [0:15];
reg [0:31] rom_O [0:15];
reg [0:31] rom_P [0:15];
reg [0:31] rom_Q [0:15];
reg [0:31] rom_R [0:15];
reg [0:31] rom_S [0:15];
reg [0:31] rom_T [0:15];
reg [0:31] rom_U [0:15];
reg [0:31] rom_V [0:15];
reg [0:31] rom_W [0:15];
reg [0:31] rom_X [0:15];
reg [0:31] rom_Y [0:15];
reg [0:31] rom_Z [0:15];
reg [0:31] rom_white [0:15];


parameter data_A = {

	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000001000000000000000000000,
	32'b00000000010100000000000000000000,
	32'b00000000100010000000000000000000,
	32'b00000001000001000000000000000000,
	32'b00000010000000100000000000000000,
	32'b00000100000000010000000000000000,
	32'b00001111111111111000000000000000,
	32'b00010000000000000100000000000000,
	32'b00100000000000000010000000000000,
	32'b01000000000000000001000000000000,
	32'b10000000000000000000100000000000
	
	};
	
	parameter data_B = {

	32'b00000001111110000000000000000000,
	32'b00000001000001000000000000000000,
	32'b00000001000000100000000000000000,
	32'b00000001000000100000000000000000,
	32'b00000001000000100000000000000000,
	32'b00000001000000100000000000000000,
	32'b00000001000001000000000000000000,
	32'b00000001111110000000000000000000,
	32'b00000001000001000000000000000000,
	32'b00000001000000100000000000000000,
	32'b00000001000000100000000000000000,
	32'b00000001000000100000000000000000,
	32'b00000001000000100000000000000000,
	32'b00000001000000100000000000000000,
	32'b00000001000001000000000000000000,
	32'b00000001111110000000000000000000
	
	};
	
	parameter data_C = {

	32'b00000000000000000000000000000000,
	32'b00000000000000010000000000000000,
	32'b00000000000000100000000000000000,
	32'b00000000000001000000000000000000,
	32'b00000000000010000000000000000000,
	32'b00000000000100000000000000000000,
	32'b00000000001000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000100000000000000000000000,
	32'b00000000100000000000000000000000,
	32'b00000000100000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000001000000000000000000000,
	32'b00000000000100000000000000000000,
	32'b00000000000010000000000000000000,
	32'b00000000000001000000000000000000
	
	};
	
	parameter data_D = {

	32'b11111110000000000000000000000000,
	32'b01000001000000000000000000000000,
	32'b01000000100000000000000000000000,
	32'b01000000010000000000000000000000,
	32'b01000000001000000000000000000000,
	32'b01000000001000000000000000000000,
	32'b01000000001000000000000000000000,
	32'b01000000001000000000000000000000,
	32'b01000000001000000000000000000000,
	32'b01000000001000000000000000000000,
	32'b01000000001000000000000000000000,
	32'b01000000001000000000000000000000,
	32'b01000000010000000000000000000000,
	32'b01000000100000000000000000000000,
	32'b01000001000000000000000000000000,
	32'b01111110000000000000000000000000
	
	};
	
	parameter data_E = {

	32'b00000000011111111110000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000011111111110000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000011111111110000000000000
	
	};
	
	parameter data_F = {

	32'b00000000011111111110000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000011111111110000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000
	
	};
	
	parameter data_G = {

	32'b00000000000000000000000000000000,
	32'b00000000000000010000000000000000,
	32'b00000000000000100000000000000000,
	32'b00000000000001000000000000000000,
	32'b00000000000010000000000000000000,
	32'b00000000000100000000000000000000,
	32'b00000000001000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000100000011111111000000000,
	32'b00000000100000000001000000000000,
	32'b00000000100000000010000000000000,
	32'b00000000010000000100000000000000,
	32'b00000000001111111000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000
	
	};
	
	parameter data_H = {

	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000011111111110000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000
	
	};
	
	parameter data_I = {

	32'b00000111111111000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000111111111100000000000000000
	
	};
	
	parameter data_J = {

	32'b00000111111100000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b01000000010000000000000000000000,
	32'b01000000100000000000000000000000,
	32'b00010001000000000000000000000000,
	32'b00001100000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000
	
	};
	
	parameter data_K = {

	32'b00000000010000000100000000000000,
	32'b00000000010000001000000000000000,
	32'b00000000010000010000000000000000,
	32'b00000000010000100000000000000000,
	32'b00000000010001000000000000000000,
	32'b00000000010010000000000000000000,
	32'b00000000010100000000000000000000,
	32'b00000000011000000000000000000000,
	32'b00000000010100000000000000000000,
	32'b00000000010010000000000000000000,
	32'b00000000010001000000000000000000,
	32'b00000000010000100000000000000000,
	32'b00000000010000010000000000000000,
	32'b00000000010000001000000000000000,
	32'b00000000010000000100000000000000,
	32'b00000000010000000010000000000000
	
	};
	
	parameter data_L = {

	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000100000000,
	32'b00000000011111111111111100000000
	
	};
	
	parameter data_M = {

	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000011000000110000000000000,
	32'b00000000010100001010000000000000,
	32'b00000000010010010010000000000000,
	32'b00000000010001000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000
	
	};
	
	parameter data_N = {

	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000011000000010000000000000,
	32'b00000000010100000010000000000000,
	32'b00000000010010000010000000000000,
	32'b00000000010001000010000000000000,
	32'b00000000010000100010000000000000,
	32'b00000000010000010010000000000000,
	32'b00000000010000001010000000000000,
	32'b00000000010000000110000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000
	
	};
	
	parameter data_O = {

	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000001100000000000000000,
	32'b00000000000010010000000000000000,
	32'b00000000001000001000000000000000,
	32'b00000000100000000010000000000000,
	32'b00000000100000000000100000000000,
	32'b00000000100000000000010000000000,
	32'b00000000001000000000100000000000,
	32'b00000000000010000010000000000000,
	32'b00000000000001111000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000
	
	};
	
	parameter data_P = {

	32'b00000001111110000000000000000000,
	32'b00000001000001000000000000000000,
	32'b00000001000000100000000000000000,
	32'b00000001000000100000000000000000,
	32'b00000001000000100000000000000000,
	32'b00000001000000100000000000000000,
	32'b00000001000001000000000000000000,
	32'b00000001111110000000000000000000,
	32'b00000001000000000000000000000000,
	32'b00000001000000000000000000000000,
	32'b00000001000000000000000000000000,
	32'b00000001000000000000000000000000,
	32'b00000001000000000000000000000000,
	32'b00000001000000000000000000000000,
	32'b00000001000000000000000000000000,
	32'b00000001000000000000000000000000
	
	};
	
	parameter data_Q = {

	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000001100000000000000000,
	32'b00000000000010010000000000000000,
	32'b00000000001000001000000000000000,
	32'b00000000100000000010000000000000,
	32'b00000000100000000000100000000000,
	32'b00000000100000000000010000000000,
	32'b00000000001000000000100000000000,
	32'b00000000000010000010000000000000,
	32'b00000000000111111111100000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000
	
	};
	
	parameter data_R = {

	32'b00000001111110000000000000000000,
	32'b00000001000001000000000000000000,
	32'b00000001000000100000000000000000,
	32'b00000001000000100000000000000000,
	32'b00000001000000100000000000000000,
	32'b00000001000000100000000000000000,
	32'b00000001000001000000000000000000,
	32'b00000001111110000000000000000000,
	32'b00000001000001000000000000000000,
	32'b00000001000000100000000000000000,
	32'b00000001000000010000000000000000,
	32'b00000001000000001000000000000000,
	32'b00000001000000000100000000000000,
	32'b00000001000000000010000000000000,
	32'b00000001000000000001000000000000,
	32'b00000001000000000000100000000000
	
	};
	
	parameter data_S = {

	32'b00000000000000000000000000000000,
	32'b00000000001111111100000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000001000000000000000000000,
	32'b00000000000100000000000000000000,
	32'b00000000000001111100000000000000,
	32'b00000000000000000100000000000000,
	32'b00000000000000000100000000000000,
	32'b00000000000000000100000000000000,
	32'b00000000000000001000000000000000,
	32'b0000000010000010000000000000000,
	32'b00000000011111100000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000
	
	};
	
	parameter data_T = {

	32'b01111111111111111100000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000000000000000000000000000000
	
	};
	
	parameter data_U = {

	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000011111111110000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000
	
	};
	
	parameter data_V = {

	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00001000000000000000100000000000,
	32'b00000100000000000001000000000000,
	32'b00000010000000000010000000000000,
	32'b00000001000000000100000000000000,
	32'b00000000100000001000000000000000,
	32'b00000000010000010000000000000000,
	32'b00000000001000100000000000000000,
	32'b00000000000101000000000000000000,
	32'b00000000000010000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000
	
	};
	
	parameter data_W = {

	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010000000010000000000000,
	32'b00000000010001000010000000000000,
	32'b00000000010010100010000000000000,
	32'b00000000010100010010000000000000,
	32'b00000000010000001110000000000000
	
	};
	
	parameter data_X = {

	32'b10000000000000010000000000000000,
	32'b01000000000000100000000000000000,
	32'b00100000000001000000000000000000,
	32'b00010000000010000000000000000000,
	32'b00001000000100000000000000000000,
	32'b00000100001000000000000000000000,
	32'b00000010010000000000000000000000,
	32'b00000001100000000000000000000000,
	32'b00000001100000000000000000000000,
	32'b00000010010000000000000000000000,
	32'b00000100001000000000000000000000,
	32'b00001000000100000000000000000000,
	32'b00010000000010000000000000000000,
	32'b00100000000001000000000000000000,
	32'b01000000000000100000000000000000,
	32'b10000000000000010000000000000000
	
	};
	
	parameter data_Y = {

	32'b10000000000000010000000000000000,
	32'b01000000000000100000000000000000,
	32'b00100000000001000000000000000000,
	32'b00010000000010000000000000000000,
	32'b00001000000100000000000000000000,
	32'b00000100001000000000000000000000,
	32'b00000010010000000000000000000000,
	32'b00000001100000000000000000000000,
	32'b00000001000000000000000000000000,
	32'b00000010000000000000000000000000,
	32'b00000100000000000000000000000000,
	32'b00001000000000000000000000000000,
	32'b00010000000000000000000000000000,
	32'b00100000000000000000000000000000,
	32'b01000000000000000000000000000000,
	32'b10000000000000000000000000000000
	
	};
	
	parameter data_Z = {

	32'b00001111111111111111111100000000,
	32'b00000000000000000000001000000000,
	32'b00000000000000000000010000000000,
	32'b00000000000000000000100000000000,
	32'b00000000000000000100000000000000,
	32'b00000000000000010000000000000000,
	32'b00000000000001000000000000000000,
	32'b00000000000100000000000000000000,
	32'b00000000010000000000000000000000,
	32'b00000001000000000000000000000000,
	32'b00000100000000000000000000000000,
	32'b00001111111111111111111100000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000
	
	};
	
	
	parameter data_white = {

	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111,
	32'b11111111111111111111111111111111
	
	};
	
	
	integer i;
	
	initial
		begin
			for (i = 0; i < 16; i = i + 1)
				begin
					rom_A [i] = data_A[(511-32*i)-:32];
					rom_B [i] = data_B[(511-32*i)-:32];
					rom_C [i] = data_C[(511-32*i)-:32];
					rom_D [i] = data_D[(511-32*i)-:32];
					rom_E [i] = data_E[(511-32*i)-:32];
					rom_F [i] = data_F[(511-32*i)-:32];
					rom_G [i] = data_G[(511-32*i)-:32];
					rom_H [i] = data_H[(511-32*i)-:32];
					rom_I [i] = data_I[(511-32*i)-:32];
					rom_J [i] = data_J[(511-32*i)-:32];
					rom_K [i] = data_K[(511-32*i)-:32];
					rom_L [i] = data_L[(511-32*i)-:32];
					rom_M [i] = data_M[(511-32*i)-:32];
					rom_N [i] = data_N[(511-32*i)-:32];
					rom_O [i] = data_O[(511-32*i)-:32];
					rom_P [i] = data_P[(511-32*i)-:32];
					rom_Q [i] = data_Q[(511-32*i)-:32];
					rom_R [i] = data_R[(511-32*i)-:32];
					rom_S [i] = data_S[(511-32*i)-:32];
					rom_T [i] = data_T[(511-32*i)-:32];
					rom_U [i] = data_U[(511-32*i)-:32];
					rom_V [i] = data_V[(511-32*i)-:32];
					rom_W [i] = data_W[(511-32*i)-:32];
					rom_X [i] = data_X[(511-32*i)-:32];
					rom_Y [i] = data_Y[(511-32*i)-:32];
					rom_Z [i] = data_Z[(511-32*i)-:32];
					rom_white [i] = data_white[(511-32*i)-:32];					
				end
		end
	
	
	always @(key_code or addr)
		begin
			case (key_code)

				8'h1c:  M  =  rom_A[addr];  //  A 
				8'h32:  M  =  rom_B[addr];  //  B 
				8'h21:  M  =  rom_C[addr];  //  C 
				8'h23:  M  =  rom_D[addr];  //  D 
				8'h24:  M  =  rom_E[addr];  //  E 
				8'h2b:  M  =  rom_F[addr];  //  F 
				8'h34:  M  =  rom_G[addr];  //  G 
				8'h33:  M  =  rom_H[addr];  //  H 
				8'h43:  M  =  rom_I[addr];  //  I 
				8'h3b:  M  =  rom_J[addr];  //  J 
				8'h42:  M  =  rom_K[addr];  //  K 
				8'h4b:  M  =  rom_L[addr];  //  L 
				8'h3a:  M  =  rom_M[addr];  //  M 
				8'h31:  M  =  rom_N[addr];  //  N 
				8'h44:  M  =  rom_O[addr];  //  O 
				8'h4d:  M  =  rom_P[addr];  //  P 
				8'h15:  M  =  rom_Q[addr];  //  Q 
				8'h2d:  M  =  rom_R[addr];  //  R 
				8'h1b:  M  =  rom_S[addr];  //  S 
				8'h2c:  M  =  rom_T[addr];  //  T 
				8'h3c:  M  =  rom_U[addr];  //  U 
				8'h2a:  M  =  rom_V[addr];  //  V 
				8'h1d:  M  =  rom_W[addr];  //  W 
				8'h22:  M  =  rom_X[addr];  //  X 
				8'h35:  M  =  rom_Y[addr];  //  Y 
				8'h1a:  M  =  rom_Z[addr];  //  Z 
	
				default:M  =  rom_white[addr];
			endcase
		end
	

endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:				Iqra University 
// Engineer: 			Kashif Inayat
// 
// Create Date:    		19-Jan-2011 
// Design Name: 
// Module Name:    		top_level 
// Project Name: 
// Target Devices:		Digilent Nexsys 2 board 
// Tool versions: 
// Description: 			This module instantiates "counter_pushbutton.v"
//								"seven_segments.v", program memory ("PM_inst") and 
//								implements a 2 to 1 multiplexer
//								"counter_pushbutton.v" outputs a counter value (9 bit) and 
//								this counter value acts as an address for program 
//								memory. The program memory can be edited here in verilog
//								code. The multiplexer selects whether counter value
//								or corresponding program memory data (instruction)
//								is diplayed on 7 segment display
//
//								INPUTS
//								-- clk- 50MHz clock from Nexsys 2 board (see ucf file)
// 							-- rst- Resets the counter to zero on low to high transition (see ucf file for pin connection)
//								-- push_button-  Increments counter on low to high transition
//								-- sel_pc- if 0, pc is displayed on 7 segment display
//												if 1, instruction (program memory data) is displayed
//												on 7 segment display.
//								
//								OUTPUTS
//								-- seven_segment- For displaying on 7 segment display
//								-- dp- For displaying on 7 segment display
//								-- an- For displaying on 7 segment display
//								
//								All outputs are for seven segment display.
//
//								For pin connections of inputs and outputs of 
//								"top_level.v" see "top_level.ucf"
//
// Dependencies: 			"counter_pushbutton.v"   "seven_segments.v"  "top_level.ucf"
//							 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module top_level(
	input clk,
	input rst,
	input push_button,
	input sel_pc,
	output [6:0] seven_segment,
	output dp,
	output [3:0] an
    );

	wire [8:0] pc;
	wire [31:0] instruction;  // contains program memory data corresponding to address "pc"
	reg [15:0] word2display;


	// instantiation of counter module

	counter_pushbutton counter_pushbutton_inst(
	.clk(clk),
	.rst(rst),
	.push_button(push_button),
	.pc(pc)
    );

	// instantiation of display module
	
	seven_segments seven_segments_inst(
	.clk(clk),
	.word2display(word2display),
	.seven_segment(seven_segment),
	.dp(dp),
	.an(an)
    );

	// Implementation of mux

	always @(*)
		begin
			if (sel_pc == 1'b0)
				word2display = {7'd0,pc};
			else
				word2display = instruction[15:0];
		end



	/////////////////////////////////////////////////////////////////////////
	// 512 x 32 program memory (512 memory location each 32 bit wide)
	// Because our single instruction is 32 bit wide 
	
	
   RAMB16_S36 #(
      .INIT(36'h000000000),  // Value of output RAM registers at startup
      .SRVAL(36'h000000000), // Output value upon SSR assertion
      .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The following INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 127
      .INIT_00(256'h00000000_00000000_00000000_20c00002_28040002_00820000_20400001_20000000),
      .INIT_01(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_02(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_03(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_04(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_05(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_06(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_07(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_08(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_09(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      // Address 128 to 255
      .INIT_10(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_11(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_12(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_13(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_14(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_15(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_16(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_17(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_18(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_19(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      // Address 256 to 383
      .INIT_20(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_21(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_22(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_23(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_24(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_25(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_26(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_27(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_28(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_29(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      // Address 384 to 511
      .INIT_30(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_31(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_32(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_33(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_34(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_35(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_36(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_37(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_38(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_39(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),

      // The next set of INITP_xx are for the parity bits
      // Address 0 to 127
      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 128 to 255
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 256 to 383
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 384 to 511
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) PM_inst (
      .DO(instruction),      	// 32-bit Data Output
      .DOP(),    					// 4-bit parity Output
      .ADDR(pc),  				// 9-bit Address Input
      .CLK(clk),    				// Clock
      .DI(),      				// 32-bit Data Input
      .DIP(),    					// 4-bit parity Input
      .EN(1'b1),      			// RAM Enable Input
      .SSR(1'b0),    			// Synchronous Set/Reset Input
      .WE(4'b0000)       		// Write Enable Input
   );

   // End of PM_inst instantiation
							
							
endmodule
